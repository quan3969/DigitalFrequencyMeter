/*************************** 数据选择 **************************/
/* 输入：	Q1			计数器1计数结果
/*     	Q2			计数器2计数结果
/*			Q3			计数器3计数结果
/*			Q4			计数器4计数结果
/*			SEL		选择输出的结果：
/*							计数器1结果（K1,K2不按）
/*							计数器2结果（K1按下）
/*							计数器3结果（K2按下）
/*							计数器4结果（K1,K2都按下）
/* 输出：	DATA 		处理后的结果
/***************************************************************/
module MUX (Q1, Q2, Q3, Q4, SEL, DATA);
	
	input [31:0] Q1, Q2, Q3, Q4;
	input [1:0] SEL;
	output DATA[31:0];
	reg [31:0] DATA;
	
	always@(SEL)
	case(SEL)
		3 : DATA <= Q1;
		1 : DATA <= Q2;
		2 : DATA <= Q3;
		0 : DATA <= Q4;
		default : DATA <= 0;
	endcase

endmodule
